
* SPICE subcircuit for bq79616_subckt_002_s37.png

.SUBCKT SUBCKT_bq79616_002_s37 PWR GND J6_PIN_1 \
+ TSREF_51 NEGSV_44 LDOIN_47 NPNB_48 BAT_1 REFHP_37 \
+ AVDD_38 CVDD_45 DVDD_49 \
+ VC0_35 VC1_33 VC2_31 VC3_29 VC4_27 VC5_25 VC6_23 VC7_21 VC8_19 VC9_17 VC10_15 VC11_13 VC12_11 VC13_9 VC14_7 VC15_5 VC16_3 \
+ CB0_34 CB1_32 CB2_30 CB3_28 CB4_26 CB5_24 CB6_22 CB7_20 CB8_18 CB9_16 CB10_14 CB11_12 CB12_10 CB13_8 CB14_6 CB15_4 CB16_2 \
+ GPIO1_61 GPIO2_60 GPIO3_59 GPIO4_58 GPIO5_57 GPIO6_56 GPIO7_55 GPIO8_54 \
+ COMHP_43 COMHN_42 COMLP_40 COMLN_41 \
+ RX_52 TX_53 NFAULT_62 \
+ BBP_64 BBN_63

* Internal Net Definitions
.NET PWR_R5_OUT
.NET LED_ANODE


* Components
R5 PWR PWR_R5_OUT 30.0

C2 TSREF_51 GND 1uF
C3 NEGSV_44 GND 0.1uF
C59 LDOIN_47 GND 0.1uF
C5 PWR_R5_OUT GND 10nF
C6 AVDD_38 GND 1uF
C7 CVDD_45 GND 4.7uF
C8 DVDD_49 GND 1uF
C9 REFHP_37 GND 1uF

R121 PWR_R5_OUT LED_ANODE 1.0k
D1 LED_ANODE J6_PIN_1 D_LED_GREEN * Assuming a generic green LED model

* Connector J6
* J6_PIN_1 is an external port connected to D1 cathode.
* Pin 2 of J6 is connected to GND directly within this subcircuit.

* IC Stub Instantiation for U1: BQ79616PAPQ1
XU1_BQ79616_stub \
+ BAT_1 CB16_2 VC16_3 CB15_4 VC15_5 CB14_6 VC14_7 CB13_8 VC13_9 CB12_10 VC12_11 CB11_12 CB10_14 VC10_15 CB9_16 VC9_17 \
+ CB8_18 VC8_19 CB7_20 VC7_21 CB6_22 VC6_23 CB5_24 VC5_25 CB4_26 VC4_27 CB3_28 VC3_29 CB2_30 VC2_31 CB1_32 VC1_33 CB0_34 VC0_35 \
+ REFHM_36 AVDD_38 AVSS_39 COMLP_40 COMLN_41 COMHN_42 COMHP_43 NEGSV_44 CVDD_45 CVSS_46 LDOIN_47 NPNB_48 DVDD_49 DVSS_50 \
+ TSREF_51 RX_52 TX_53 GPIO8_54 GPIO7_55 GPIO6_56 GPIO5_57 GPIO4_58 GPIO3_59 GPIO2_60 GPIO1_61 NFAULT_62 BBN_63 BBP_64 PAD_65 \
+ BQ79616_stub

.ENDS SUBCKT_bq79616_002_s37

* Stub subcircuit for U1 (BQ79616PAPQ1)
* Internal behavior intentionally omitted; to be filled by another agent.
.SUBCKT BQ79616_stub \
+ BAT_1 CB16_2 VC16_3 CB15_4 VC15_5 CB14_6 VC14_7 CB13_8 VC13_9 CB12_10 VC12_11 CB11_12 CB10_14 VC10_15 CB9_16 VC9_17 \
+ CB8_18 VC8_19 CB7_20 VC7_21 CB6_22 VC6_23 CB5_24 VC5_25 CB4_26 VC4_27 CB3_28 VC3_29 CB2_30 VC2_31 CB1_32 VC1_33 CB0_34 VC0_35 \
+ REFHM_36 AVDD_38 AVSS_39 COMLP_40 COMLN_41 COMHN_42 COMHP_43 NEGSV_44 CVDD_45 CVSS_46 LDOIN_47 NPNB_48 DVDD_49 DVSS_50 \
+ TSREF_51 RX_52 TX_53 GPIO8_54 GPIO7_55 GPIO6_56 GPIO5_57 GPIO4_58 GPIO3_59 GPIO2_60 GPIO1_61 NFAULT_62 BBN_63 BBP_64 PAD_65

* Connect the U1 pins that are tied to ground in this schematic directly to GND.
* This implies these pins are internal to the U1 model stub, but connected to the parent\'s GND.
R_PAD_65_GND PAD_65 GND 0 * Assuming a 0 Ohm connection to the main subcircuit\'s GND
R_REFHM_36_GND REFHM_36 GND 0
R_AVSS_39_GND AVSS_39 GND 0
R_CVSS_46_GND CVSS_46 GND 0
R_DVSS_50_GND DVSS_50 GND 0

.ENDS BQ79616_stub

* Generic diode model for D1
.MODEL D_LED_GREEN D
